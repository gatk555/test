Verilog-controlled simple timer.

* This sub-circuit simulates the NE555 timer IC, with the digital part
* as a GHDL entity.

.subckt NE555 trigger threshold reset control output discharge vcc ground

* Resistor chain

r1 vcc control 5k
r2 control trigger_ref 5k
r3 trigger_ref ground 5k

* Two XSPICE ADC instances serve as comparators.

.model comparator adc_bridge(in_low = -0.0001 in_high = 0.0001)
athresh_comparator [%vd threshold control] [over_threshold] comparator
atrigger_comparator [%vd trigger_ref trigger] [under_trigger] comparator

* A tiny VHDL module supplies the flip-flop.

adut [ under_trigger over_threshold reset ] [ output qbar ] logic
.model logic d_cosim simulation="timer_core" sim_args=["555"]

* The discharge transistor and its base resistor.

rbase qbar discharge_base 10k
qdischarge discharge discharge_base ground npn_transistor
.model npn_transistor npn

.ends ; Ends subcircuit NE555


* The usual 555 oscillator with threshold connected to discharge.

.param vcc=12

X555 trigger_threshold trigger_threshold reset control output discharge vcc 0 ne555

r1 vcc discharge 10k
r2 discharge trigger_threshold 10k
Ct trigger_threshold 0 1uF ic=0

* A resistive load forces analog output.

rload output 0 1k

* A voltage source for power.

Vcc vcc 0 {vcc}

* Pulse the Reset signal low for 2uS each 51mS

Vpulse reset 0 PULSE {vcc} 0.2 0 1u 1u 2u 51m

.tran 10u 200m uic
.control
iplot -d 200 trigger_threshold output
*run
.endc
.end
