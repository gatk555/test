Test divide by 3 VHDL code

adut null [clk cout] d3
.model d3 d_cosim simulation=./wrapper.so

r1 clk 0 29k
r2 cout 0 29k

.tran 100n 10u
.control
*run
*plot clk cout+1.5
.endc
.end

